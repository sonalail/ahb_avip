`ifndef AHBENVIRONMENTPACKAGE_INCLUDED_
`define AHBENVIRONMENTPACKAGE_INCLUDED_

package AhbEnvironmentPackage;
  
  import AhbGlobalPackage::*;
  import AhbMasterPackage::*;
  import AhbSlavePackage::*;

  `include "AhbVirtualSequencer.sv"
  `include "AhbScoreboard.sv"
  `include "AhbEnvironment.sv"

endpackage : AhbEnvironmentPackage

`endif
