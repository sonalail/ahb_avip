

`ifndef AHBMASTERPACKAGE_INCLUDED_
`define AHBMASTERPACKAGE_INCLUDED_

package AhbMasterPackage;

  `include "uvm_macros.svh"

  import uvm_pkg::*;
  import AhbGlobalPackage::*;

  `include "AhbMasterAgentConfig.sv"
  `include "AhbMasterTransaction.sv"
  `include "AhbMasterSequenceItemConverter.sv"
  `include "AhbMasterConfigConverter.sv"
  `include "AhbMasterSequencer.sv"
  `include "AhbMasterDriverProxy.sv"
  `include "AhbMasterMonitorProxy.sv"
  `include "AhbMasterCoverage.sv"
  `include "AhbMasterAgent.sv"
  
endpackage : AhbMasterPackage

`endif


