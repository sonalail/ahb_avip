`ifndef AHBBASETESTPACKAGE_INCLUDED_
`define AHBBASETESTPACKAGE_INCLUDED_

package AhbBaseTestPackage;

  `include "uvm_macros.svh"
  import uvm_pkg::*;

  import AhbGlobalPackage::*;
  import AhbMasterPackage::*;
  import AhbSlavePackage::*; 
  import AhbEnvironmentPackage::*;
  import AhbMasterSequencePackage::*;
  import AhbSlaveSequencePackage::*;
  import AhbVirtualSequencePackage::*;

  `include "AhbBaseTest.sv"
  `include "AhbWriteTest.sv"
  `include "AhbReadTest.sv"
  `include "AhbSingleWriteTest.sv"
  `include "AhbSingleReadTest.sv"
  `include "AhbWriteWithBusyTest.sv"
  `include "AhbReadWithBusyTest.sv"


endpackage : AhbBaseTestPackage

`endif
