`ifndef HVLTOP_INCLUDED_
`define HVLTOP_INCLUDED_

module HvlTop;

  import AhbBaseTestPackage::*;
  
    run_test("AhbBaseTest");
  end

endmodule : HvlTop

`endif
